module multiplier(a, b, z);
    input [2:0] a;
    input [2:0] b;
    output reg [5:0] z;

    always @(a, b) begin
        case ({a, b})
            6'b000000: z <= 6'b000000; // 0 * 0 = 0
            6'b000001: z <= 6'b000000; // 0 * 1 = 0
            6'b000010: z <= 6'b000000; // 0 * 2 = 0
            6'b000011: z <= 6'b000000; // 0 * 3 = 0
            6'b000100: z <= 6'b000000; // 0 * 4 = 0
            6'b000101: z <= 6'b000000; // 0 * 5 = 0
            6'b000110: z <= 6'b000000; // 0 * 6 = 0
            6'b000111: z <= 6'b000000; // 0 * 7 = 0
            6'b001000: z <= 6'b000000; // 1 * 0 = 0
            6'b001001: z <= 6'b000001; // 1 * 1 = 1
            6'b001010: z <= 6'b000010; // 1 * 2 = 2
            6'b001011: z <= 6'b000011; // 1 * 3 = 3
            6'b001100: z <= 6'b000100; // 1 * 4 = 4
            6'b001101: z <= 6'b000101; // 1 * 5 = 5
            6'b001110: z <= 6'b000110; // 1 * 6 = 6
            6'b001111: z <= 6'b000111; // 1 * 7 = 7
            6'b010000: z <= 6'b000000; // 2 * 0 = 0
            6'b010001: z <= 6'b000010; // 2 * 1 = 2
            6'b010010: z <= 6'b000100; // 2 * 2 = 4
            6'b010011: z <= 6'b000110; // 2 * 3 = 6
            6'b010100: z <= 6'b001000; // 2 * 4 = 8
            6'b010101: z <= 6'b001010; // 2 * 5 = 10
            6'b010110: z <= 6'b001100; // 2 * 6 = 12
            6'b010111: z <= 6'b001110; // 2 * 7 = 14
            6'b011000: z <= 6'b000000; // 3 * 0 = 0
            6'b011001: z <= 6'b000011; // 3 * 1 = 3
            6'b011010: z <= 6'b000110; // 3 * 2 = 6
            6'b011011: z <= 6'b001001; // 3 * 3 = 9
            6'b011100: z <= 6'b001100; // 3 * 4 = 12
            6'b011101: z <= 6'b001111; // 3 * 5 = 15
            6'b011110: z <= 6'b010010; // 3 * 6 = 18
            6'b011111: z <= 6'b010101; // 3 * 7 = 21
            6'b100000: z <= 6'b000000; // 4 * 0 = 0
            6'b100001: z <= 6'b000100; // 4 * 1 = 4
            6'b100010: z <= 6'b001000; // 4 * 2 = 8
            6'b100011: z <= 6'b001100; // 4 * 3 = 12
            6'b100100: z <= 6'b010000; // 4 * 4 = 16
            6'b100101: z <= 6'b010100; // 4 * 5 = 20
            6'b100110: z <= 6'b011000; // 4 * 6 = 24
            6'b100111: z <= 6'b011100; // 4 * 7 = 28
            6'b101000: z <= 6'b000000; // 5 * 0 = 0
            6'b101001: z <= 6'b000101; // 5 * 1 = 5
            6'b101010: z <= 6'b001010; // 5 * 2 = 10
            6'b101011: z <= 6'b001111; // 5 * 3 = 15
            6'b101100: z <= 6'b010100; // 5 * 4 = 20
            6'b101101: z <= 6'b011001; // 5 * 5 = 25
            6'b101110: z <= 6'b011110; // 5 * 6 = 30
            6'b101111: z <= 6'b100011; // 5 * 7 = 35
            6'b110000: z <= 6'b000000; // 6 * 0 = 0
            6'b110001: z <= 6'b000110; // 6 * 1 = 6
            6'b110010: z <= 6'b001100; // 6 * 2 = 12
            6'b110011: z <= 6'b010010; // 6 * 3 = 18
            6'b110100: z <= 6'b011000; // 6 * 4 = 24
            6'b110101: z <= 6'b011110; // 6 * 5 = 30
            6'b110110: z <= 6'b100100; // 6 * 6 = 36
            6'b110111: z <= 6'b101010; // 6 * 7 = 42
            6'b111000: z <= 6'b000000; // 7 * 0 = 0
            6'b111001: z <= 6'b000111; // 7 * 1 = 7
            6'b111010: z <= 6'b001110; // 7 * 2 = 14
            6'b111011: z <= 6'b010101; // 7 * 3 = 21
            6'b111100: z <= 6'b011100; // 7 * 4 = 28
            6'b111101: z <= 6'b100011; // 7 * 5 = 35
            6'b111110: z <= 6'b101010; // 7 * 6 = 42
            6'b111111: z <= 6'b110001; // 7 * 7 = 49
            default: z <= 0;
        endcase
    end
endmodule
